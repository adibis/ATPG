1 1 0 2 0
1 2 0 1 0
1 3 0 1 0
1 4 0 1 0
2 5 1 1 
2 6 1 1
0 7 2 2 3 2 3 4 
2 8 1 7
2 9 1 7
0 10 4 2 2 6 8
0 11 5 1 1 9 
2 12 1 10
2 13 1 10
3 14 6 0 2 5 12 
3 15 2 0 2 11 13
