1 1 0 2 0
1 2 0 2 0
2 4 1 1
2 5 1 1
2 6 1 2
2 7 1 2
2 8 1 3
2 9 1 3
3 10 2 0 3 4 6 8
1 3 0 2 0
3 11 2 0 3 5 7 9
