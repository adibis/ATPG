1 1  0 1  0
1 2  0 1  0
1 3  0 2  0
2 4  1 3
2 5  1 3
1 6  0 1  0
1 7  0 2  0
2 8  1 7
2 9  1 7
1 10 0 1  0
1 11 0 1  0
1 12 0 1  0
0 13 6 1  3 1 2 4
0 14 6 1  3 5 6 8
0 15 6 2  3 9 10 11
2 16 1 15
2 17 1 15
0 18 6 1  3 13 14 16
0 19 3 1  2 17 12
3 20 2 0  2 18 19
