1 1 0 1 0
1 2 0 1 0
1 3 0 1 0
1 4 0 1 0
1 5 0 2 0
2 6 1 5
2 7 1 5
0 8 3 1 2 1 2
0 9 7 1 2 4 6
0 10 3 2 2 3 9
2 11 1 10
2 12 1 10
0 13 5 1 1 11
0 14 2 1 3 12 7 17
0 15 3 1 2 8 13
3 16 6 0 2 15 14
1 17 0 1 0